*****************************************************************************************
* Library Name: subADAC
* Cell Name: subADC
* View Name: schematic
*****************************************************************************************

.SUBCKT subADC vref vIref clk vddl vssl vip out1 out2 out3 out4 out5 out6

IIin vddl Iin 2u

* 分压电路
R1 pot1 vIref 300k
R2 pot2 pot1 200k
R3 pot3 pot2 200k
R4 pot4 pot3 200k
R5 pot5 pot4 200k
R6 pot6 pot5 200k
R7 vref pot6 300k
*R8 vref pot7 5k

* 比较电路
xc1 Iin clk vssl out1 vddl pot1 vip comparator_preamp $-1.0V
xc2 Iin clk vssl out2 vddl pot2 vip comparator_preamp $-0.6V
xc3 Iin clk vssl out3 vddl pot3 vip comparator_preamp $-0.2V
xc4 Iin clk vssl out4 vddl pot4 vip comparator_preamp $0.2V
xc5 Iin clk vssl out5 vddl pot5 vip comparator_preamp $0.6V
xc6 Iin clk vssl out6 vddl pot6 vip comparator_preamp $1.0V

$ 滤波电路
c11 pot1 0 10u
c12 pot2 0 10u
c13 pot3 0 10u
c14 pot4 0 10u
c15 pot5 0 10u
c16 pot6 0 10u

c21 out1 0 10p
c22 out2 0 10p
c23 out3 0 10p
c24 out4 0 10p
c25 out5 0 10p
c26 out6 0 10p

.ENDS

*****************************************************************************************
* Library Name: subADAC
* Cell Name: subDAC
* View Name: schematic
*****************************************************************************************

.SUBCKT subDACa vdd vss vin out1 out2 out3 out4 out5 out6 out

xI Vp Vn Ivin vdd vss / OPAMP
R1 Vn vin 1M
R2 Vn Ivin 1M
R3 Vp 0 10k

Ra out1 in1 1M
Rb out2 in1 1M
Rc out3 in1 1M
Rd out4 in1 1M
Re out5 in1 1M
Rf out6 in1 1M
Ri Ivin in1 62k

XI1 0 in1 outm vdd vss / OPAMP
XI2 outm in2 out vdd vss / OPAMP

RA1 in1 outm 100k
RA21 out in2 150k
RA22 in2 0 100k

.ENDS

.SUBCKT subDAC vref vIref vdd vss vin out1 out2 out3 out4 out5 out6 out

*开关电路决定电源高低
xs1 vdd vss out1 vref ina / BOOSTRAP
xs2 vdd vss out2 vref inb / BOOSTRAP
xs3 vdd vss out3 vref inc / BOOSTRAP
xs4 vdd vss out4 vref ind / BOOSTRAP
xs5 vdd vss out5 vref ine / BOOSTRAP
xs6 vdd vss out6 vref inf / BOOSTRAP

R1 Vn ina 2k
R2 Vn inb 2k
R3 Vn inc 2k
R4 Vn ind 2k
R5 Vn ine 2k
R6 Vn inf 2k

Rno Vn out 1k

XI vin Vn out vdd vss / OPAMP

.ENDS

************************************************
* ��������ģ���·������                        
* ��������������ϵͳ������·��                  
************************************************
* ���������¿������ܽ�                        
************************************************
* ����������ѧ�����硡2020                      
************************************************          
*
*****************************************************************************************
* Library Name: comparator
* Cell Name: INV
* View Name: schematic
*****************************************************************************************
* CMOS inverter
.subckt INV vdda gnda  in out 
MPM2 out in vdda vdda p18 W=4u L=180n m=1
MNM1 out in gnda gnda n18 W=2u L=180n m=1
.ends

* CMOS inverter with larger delay
.subckt INV2 vdda gnda  in out 
MPM2 out in vdda vdda p18 W=20u L=900n m=1
MNM1 out in gnda gnda n18 W=10u L=900n m=1
.ends

* CMOS inverter with further larger delay based on INV2 (5x of W&L)
* 10x larger of delay
* clk1d ����� clk1���½����ӳ�Լ2.3ns
* �������INV���½����ӳ�Լ0.25ns
.subckt INV1 vdda gnda  in out 
x1 vdda gnda  in    net01 / INV2
x2 vdda gnda  net01 net02 / INV2 
x3 vdda gnda  net02 net03 / INV2
x4 vdda gnda  net03 net04 / INV2 
x5 vdda gnda  net04 net05 / INV2 
x6 vdda gnda  net05 net06 / INV2 
x7 vdda gnda  net06 out   / INV2 
.ends

* CMOS switch
.subckt SWITCHb vdda gnda  s  in out 
x1 vdda gnda  s s_inv / INV
m1 out s     in gnda n18 W=2u L=180n m=1
m2 out s_inv in vdda p18 W=4u L=180n m=1
.ends

*****************************************************************************************
* Library Name: comparator
* Cell Name: NAND
* View Name: schematic
*****************************************************************************************
* CMOS nand
.SUBCKT NAND vdda gnda  A B out
MPM2 out A vdda vdda p18 W=4u L=180n m=1
MPM1 out B vdda vdda p18 W=4u L=180n m=1
MNM1 net01 B gnda gnda n18 W=2u L=180n m=1
MNM2 out A net01 gnda n18 W=2u L=180n m=1
.ENDS

* CMOS and
.SUBCKT AND vdda gnda  A B out
x1 vdda gnda  A B  outn / NAND
x2 vdda gnda  outn out  / INV 
.ENDS

* CMOS buffer
.SUBCKT buffer vdda gnda in out
x1 vdda gnda  in  in_inv / INV
x2 vdda gnda  in_inv out / INV 
.ENDS

* non-overlap clock generation
.subckt CLOCKb vdda gnda  clkin clk1 clk1d clk2 clk2d
xa1  vdda gnda clkin net05 net01  / NAND
xa2  vdda gnda net01 net03 net04  / NAND
xa3  vdda gnda net06 net07 net08  / NAND
xa4  vdda gnda net08 net10 net11  / NAND

xi1  vdda gnda net01 net02        / INV
xi2  vdda gnda net02 net03        / INV1
xi3  vdda gnda net08 net09        / INV
xi4  vdda gnda net09 net10        / INV1
xi5  vdda gnda clk2d net05        / INV1
xi6  vdda gnda clk1d net06        / INV1
xi7  vdda gnda clkin net07        / INV

xb1  vdda gnda net02 clk1         / BUFFER  
xb2  vdda gnda net04 clk1d        / BUFFER  
xb3  vdda gnda net09 clk2         / BUFFER  
xb4  vdda gnda net11 clk2d        / BUFFER  
.ends
****************************
* in use
****************************
* non-overlap clock generation
.subckt CLOCKa vdda gnda  clkin clk1 clk1d clk2 clk2d
xa1  vdda gnda net12 net05 net01  / NAND
xa2  vdda gnda net01 net03 net04  / NAND
xa3  vdda gnda net06 net07 net08  / NAND
xa4  vdda gnda net08 net10 net11  / NAND

xi1  vdda gnda net01 net02        / INV
xi2  vdda gnda net02 net03        / INV1
xi3  vdda gnda net08 net09        / INV
xi4  vdda gnda net09 net10        / INV1
xi5  vdda gnda net10 net05        / INV1
xi6  vdda gnda net03 net06        / INV1
xi7  vdda gnda clkin net07        / INV
xi8  vdda gnda net07 net12        / INV

xb1  vdda gnda net02 clk1         / BUFFER  
xb2  vdda gnda net04 clk1d        / BUFFER  
xb3  vdda gnda net09 clk2         / BUFFER  
xb4  vdda gnda net11 clk2d        / BUFFER  
.ends

* latch comparator
* if vip>vin then voutp=HIGH voutn=LOW
* if vip<vin then voutp=LOW  voutn=HIGH
.SUBCKT comparator vdda gnda clk vip vin voutp voutn
xa1 vdda gnda net01  voutn voutp  / NAND
xa2 vdda gnda net02  voutp voutn  / NAND

MM1 net03 vip   gnda gnda n18 W=20u L=180n m=1
MM2 net03 net04 gnda gnda n18 W=20u L=180n m=1
MM3 net04 net03 gnda gnda n18 W=20u L=180n m=1
MM4 net04 vin   gnda gnda n18 W=20u L=180n m=1

MM5 net01 clk net03 gnda n18 W=30u L=180n m=1
MM6 net02 clk net04 gnda n18 W=30u L=180n m=1

MM7 net01 clk   vdda vdda p18 W=60u L=180n m=1
MM8 net01 net02 vdda vdda p18 W=60u L=180n m=1
MM9 net02 net01 vdda vdda p18 W=60u L=180n m=1
MM10 net02 clk  vdda vdda p18 W=60u L=180n m=1
.ENDS

*****************************************************************************************
* Library Name: comparator
* Cell Name: comparatormove
* View Name: schematic
*****************************************************************************************

.SUBCKT comparatormove clk gnda out vdda vin vip	*������̬�Ƚ�����·
XI2 vdda gnda net048 net045 / INV
XI3 vdda gnda net045 out / INV
XI0 vdda gnda outp1 net048 net049  / NAND
XI1 vdda gnda net049 outn1 net048  / NAND
MM9 outp1 outn1 vdda vdda p18 W=60u L=180n m=1
MM10 outp1 clk vdda vdda p18 W=60u L=180n m=1
MM8 outn1 outp1 vdda vdda p18 W=60u L=180n m=1
MM7 outn1 clk vdda vdda p18 W=60u L=180n m=1
MM4 net40 vin gnda gnda n18 W=20u L=180n m=1
MM3 net40 net42 gnda gnda n18 W=20u L=180n m=1
MM6 outp1 clk net40 gnda n18 W=30u L=180n m=1
MM5 outn1 clk net42 gnda n18 W=30u L=180n m=1
MM2 net42 net40 gnda gnda n18 W=20u L=180n m=1
MM1 net42 vip gnda gnda n18 W=20u L=180n m=1
.ENDS

*****************************************************************************************
* Library Name: comparator
* Cell Name: pre_amp
* View Name: schematic
*****************************************************************************************

.SUBCKT pre_amp Idc_2u gnda vdda vin vip voutn voutp //����Ԥ�Ŵ�����·
MM4 voutn voutp vdda vdda p18 W=1u L=1u m=1
MM5 voutp voutn vdda vdda p18 W=1u L=1u m=1
MM6 voutp voutp vdda vdda p18 W=1.8u L=1u m=1
MM3 voutn voutn vdda vdda p18 W=1.8u L=1u m=1
MM1 voutn vip net27 gnda n18 W=4u L=2u m=1
MM2 voutp vin net27 gnda n18 W=4u L=2u m=1
MM0 net27 Idc_2u gnda gnda n18 W=8u L=2u m=1
MMbias Idc_2u Idc_2u gnda gnda n18 W=4u L=2u m=1
.ENDS
